LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
--
--    .. hwt-autodoc::
--    
ENTITY ParametrizationExample IS
    GENERIC(
        PARAM_0 : INTEGER := 0;
        PARAM_10 : INTEGER := 10;
        PARAM_1_sll_512 : STD_LOGIC_VECTOR(512 DOWNTO 0) := "100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
        PARAM_1_sll_512_py_int : STRING := "13407807929942597099574024998205846127479365820592393377723561443721764030073546976801874298166903427690031858186486050853753882811946569946433649006084096"
    );
    PORT(
        din : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
        dout : OUT STD_LOGIC_VECTOR(19 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE rtl OF ParametrizationExample IS
BEGIN
    dout <= din & din;
    ASSERT PARAM_0 = 0 REPORT "Generated only for this value" SEVERITY failure;
    ASSERT PARAM_10 = 10 REPORT "Generated only for this value" SEVERITY failure;
    ASSERT PARAM_1_sll_512 = "100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" REPORT "Generated only for this value" SEVERITY failure;
    ASSERT PARAM_1_sll_512_py_int = "13407807929942597099574024998205846127479365820592393377723561443721764030073546976801874298166903427690031858186486050853753882811946569946433649006084096" REPORT "Generated only for this value" SEVERITY failure;
END ARCHITECTURE;
