package c is
end package;

