package body a is
end a;
