use work.b.all;

package a is 
end package;

