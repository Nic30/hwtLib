package body c is
end c;
