package body b is
end b;
