use work.c.all;

package b is
end package;

